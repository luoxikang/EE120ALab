// Verilog test fixture created from schematic B:\EE120A\Lab2Part2A\Part2A.sch - Wed Oct 09 22:22:40 2019

`timescale 1ns / 1ps

module Part2A_Part2A_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   Part2A UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
